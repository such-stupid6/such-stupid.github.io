B�Q��9G|<eUm�l�&�)��\���«p����;I�\L��0(��M*�|֨ĥ��`F�k��
]�(����.���C������$ђEd�s%�L`�����'���������L���ܬ�$�Y�H{?�T�Z���ԭqxt|xx���R<L���RGF� �� �z(�t�}q�%U�z��I�j
��3y!g��o���|�:��n��&?��Xҝ���о�A�w쐾)��N�L� �0Xs1r�Z�$t�F"MHѹ���/ۉM��Y0�H�˱��~|P�JB�%j}B�6��
��"�3�>+9�9�K�.v�B�5�f'8��uk�cWɢ&Cl�Sd�g�X@Uk&v�s3j�Js����U�E�[�*���a�� �';t��� �05��:��ϲ݉�
�۩d������\X{��T�-�;�U�i+�E���e�/�Zb2���%��{�,��Z:�+L����1ep�o�MDI@,�߯������j�;��4�f)K2c�j�nL\�,��,�#��w�v�&���c�{���w���aKr���sg���f`���n�@�9'��6\�P��v�}�K����M9t% ��A2��kb\�UQN�� �<81�=�״�l&�Y2؅��ž�}�3m;c�u�+;�5�A%��*E��!���XPAݣ�t�SZ,�C4���q�:%�W�i�NC���Sge����r>�P�d=���� s��4�dSuF�%S�׭H��jpGb(�0�ˢJ�wΘ��5u6{�4�/�&@5�BI�de�aF�FnR� �n��i�DJ%�i�fp&�����/��\�&��0���_�����{|o
��&���e���F\4R�i*�t�L4��8#�U:�ӝ�\l4sNR���ʓAܞdJj�c��S����H"�#\�����rD?G��S��*��iڻ�h�$��CM�W����鼱�6�#�O���H��
4�I��"��(~*m�1S
���4>h�����ڎj��o/&w��O�9���Mx��6��W��3�$�J�l2�)O�@\ɪ��h*�2�G*���X��Rq�N(L�y�G/0p����{ �JT^��cx��
�\!��(��#w��)}&�p��h�
������)�!�hr@���=+��O� ��Q��(�t#��V/�*�JhUtw�;���u���jQ�\F`=ㅰ�7��*o��%F�A�|�Yɤ������7�_-+��٭�;�hĶt��m5T|vI�{�b��X^��ƈ���j>�颼�$c�8���$��b��y�� v2F��4����h���!���R��:{Q�I߭b�Sz�)ȧ"�N�tͺQ���6q:���$ç;���>����\��&��P����C�K�6-�	��N�)�#�@�"U����h���)�h��Z=r�[�W���D��4��r����=%ɧ�����w&����cB\��Ig	uJ��Y+rDC5,Ҙk�Ffg������W,vj�#�Lϥ�nj&L7�;�!���d�r�2�3p�}�J>�5ܖmPXM�)�y�L�N�K����O��T�ڔ��C
�b+s�9�-�əi|S��c=��8L��!b�\(u%�aU�ݸv�z��ţ�ob�����3F��e3��1T	+!�I�3����C����a�WZ���[��H�-V�+���� �҆veۈ��ƌ����gD�3�~=�J����a�a1��ɀ�����U�������0M��<�O�H����*@?3@@���(qFה��s��?i�Yĺnkn&���{�m�r��9�x3��Mi4�N�l����pe<�<����8띏A�T&pU6\A�iL���+Y"�ҝ�?�"�l�E�n"�ƃ,J���Ƥ����ė	[P�Q��.� ΁�V�C$o���s�0:mV�84@��]��&��QDU��j�7i��?o'�5Z�Nz�o��؁F8��n�qv�D�ϸ��=P"�}4�FՃ�5��`&yi]wLL�߷J�0\��[�!]���"�+���M˹�����y'f��ş!�N^u#?A�W�0�������s��)���^�Z�܅X���w)i��w��l�����W(���Ñ�P��Xj9�RVCL�I�R�=�wω�G���D:�o�O��y~�<�9i��1M��`<%ؖڻ���a $mr�����à��.O��?��|h��Gd�='�hW��wv�f!��HR[��3̀����!f���� -9��N���)@�B���5ߺ^�I�N�Q�|�`BL�	4�~E	$W�u6��6ї����?e�&��R86�I�3_��:a� F�
��@��6�ܳ	���h#��1Z�]kt�e���a[���|լZ�f��#���W���߶;=��T���=B��z:���3� �[�Q}5�w,ឍ;��I���P%����r���<#����[�R���Lr�VS@�n$�����B<%OX�ֹ�t�K���U\ܔ��=d�7PL�����}N�<w��5O奉c�_��G��фn�o2��f�)v�$��$K_)d3uEyQ$�deO&����c��ƌ�&%�t����Tz(�&�ԸJ�cbIh�"HR)؊�Ρ�ԓ�u�6�zoEMK�8��:�������K��F�,���%Q�{��hc�~)n��X�TJ��G��L!�y�����V�&&O�����5_:��Q�������u��,7��/	7ʡ���=�,���'&�b�]&�{�&��HO����!�q����]�P�B��M���Oc�}��9'����.u�ِ4<6Q
b* A��)*��&��"�:̝ͫ���}���U�k����2�4��vh�{�%ƜnH�;�0/�5|-zC���k�?�Ƭ��Hy��zS�"�4%tð�6l��S��#PI�f)�iҴb۫���]XV��if���a��=�%k��,�VQ�-�0L�Yfؗ�s�5����_v���p�i���Czry~��0�@�}�e.��i�z/��H��e]-�u�cn��	�"���n�
o�ߛ�U�p60/���x�A����/|F����=p���2f*�	��2ӹ�1W�$�;�V�`�m��s�.���-U,an^���{�d3	��a�CFѶ��(O������N16F0F<!v1�哩����(���3X@�J��ɻ̷���H׍�ʠ��Cg��	�#JY��8�Fޛ��A�Wp0ycF�� ë"M \Cٲs�km�e����{`��踦����_�U���~��8BXJ�.�~4�<�F� x݊���^=p�ha��7P�=�d��əM�+Y�he�\�M��l&���:��O��P��|�.�5�<��÷$�3�=&�+��xJ�819�8<lqvc�f�ȱh �Ξ�;k�R£Up���7��{)拳?b<�Z�2>�I e����.��1����ĕL3��d
c�%.ϓ��x�Cc� I'SҴY	����<�ʞk�����![�w��hɧ�Oxr�kΛ����Uhz���Lٙ��Z'p:i\��&�h�[,l�3�.����rS����!y;���CF.���j�#<G��,������k�z,hB�c������uA��7���l�m�k<�zNRi������'�;ьXo!